LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LAB_EXAM1 IS
port(
SW:IN STD_LOGIC_VECTOR (7 DOWNTO 0);
LEDG:OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
LEDR:OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
);

END LAB_EXAM1;

ARCHITECTURE Behavior OF LAB_EXAM1 IS
BEGIN
LEDG<=SW;
LEDR<=SW;
END Behavior;
